module vivado_is_so_smart (
	input wire wire1_in,
	input wire wire2_in,
	output wire wire1_out,
	output wire wire2_out
);
	assign wire1_out = wire1_in;
	assign wire2_out = wire2_in;
endmodule
